//////////////////////////////////////////////////////////////////////
//          ██╗       ██████╗   ██╗  ██╗    ██████╗            		//
//          ██║       ██╔══█║   ██║  ██║    ██╔══█║            		//
//          ██║       ██████║   ███████║    ██████║            		//
//          ██║       ██╔═══╝   ██╔══██║    ██╔═══╝            		//
//          ███████╗  ██║  	  ██║  ██║    ██║  	           		//
//          ╚══════╝  ╚═╝  	  ╚═╝  ╚═╝    ╚═╝  	           		//
//                                                             		//
// 	2024 Advanced VLSI System Design, advisor: Lih-Yih, Chiou		//
//                                                             		//
//////////////////////////////////////////////////////////////////////
//                                                             		//
// 	Autor: 			TZUNG-JIN, TSAI (Leo)				  	   		//
//	Filename:		 AXI.sv			                            	//
//	Description:	Top module of AXI	 							//
// 	Version:		1.0	    								   		//
//////////////////////////////////////////////////////////////////////
// `include "AXI_define.svh"

/*
`include "WriteAddress.sv"
`include "WriteData.sv"
`include "WriteRespone.sv"
`include "ReadData.sv"
`include "ReadAddress.sv"
`include "DefaultSlave.sv"
*/

`include "../src/AXI/WriteAddress.sv"
`include "../src/AXI/WriteData.sv"
`include "../src/AXI/WriteRespone.sv"
`include "../src/AXI/ReadData.sv"
`include "../src/AXI/ReadAddress.sv"
`include "../src/AXI/DefaultSlave.sv"


module AXI(

	input ACLK,
	input ARESETn,

	//SLAVE INTERFACE FOR MASTERS
	
	//WRITE ADDRESS
	input [`AXI_ID_BITS-1:0] AWID_M1,
	input [`AXI_ADDR_BITS-1:0] AWADDR_M1,
	input [`AXI_LEN_BITS-1:0] AWLEN_M1,
	input [`AXI_SIZE_BITS-1:0] AWSIZE_M1,
	input [1:0] AWBURST_M1,
	input AWVALID_M1,
	output logic AWREADY_M1,
	
	//WRITE DATA
	input [`AXI_DATA_BITS-1:0] WDATA_M1,
	input [`AXI_STRB_BITS-1:0] WSTRB_M1,
	input WLAST_M1,
	input WVALID_M1,
	output logic WREADY_M1,
	
	//WRITE RESPONSE
	output logic [`AXI_ID_BITS-1:0] BID_M1,
	output logic [1:0] BRESP_M1,
	output logic BVALID_M1,
	input BREADY_M1,

	//READ ADDRESS0
	input [`AXI_ID_BITS-1:0] ARID_M0,
	input [`AXI_ADDR_BITS-1:0] ARADDR_M0,
	input [`AXI_LEN_BITS-1:0] ARLEN_M0,
	input [`AXI_SIZE_BITS-1:0] ARSIZE_M0,
	input [1:0] ARBURST_M0,
	input ARVALID_M0,
	output logic ARREADY_M0,
	
	//READ DATA0
	output logic [`AXI_ID_BITS-1:0] RID_M0,
	output logic [`AXI_DATA_BITS-1:0] RDATA_M0,
	output logic [1:0] RRESP_M0,
	output logic RLAST_M0,
	output logic RVALID_M0,
	input RREADY_M0,
	
	//READ ADDRESS1
	input [`AXI_ID_BITS-1:0] ARID_M1,
	input [`AXI_ADDR_BITS-1:0] ARADDR_M1,
	input [`AXI_LEN_BITS-1:0] ARLEN_M1,
	input [`AXI_SIZE_BITS-1:0] ARSIZE_M1,
	input [1:0] ARBURST_M1,
	input ARVALID_M1,
	output logic ARREADY_M1,
	
	//READ DATA1
	output logic [`AXI_ID_BITS-1:0] RID_M1,
	output logic [`AXI_DATA_BITS-1:0] RDATA_M1,
	output logic [1:0] RRESP_M1,
	output logic RLAST_M1,
	output logic RVALID_M1,
	input RREADY_M1,

	//MASTER INTERFACE FOR SLAVES
	//WRITE ADDRESS0
	output logic [`AXI_IDS_BITS-1:0] AWID_S0,
	output logic [`AXI_ADDR_BITS-1:0] AWADDR_S0,
	output logic [`AXI_LEN_BITS-1:0] AWLEN_S0,
	output logic [`AXI_SIZE_BITS-1:0] AWSIZE_S0,
	output logic [1:0] AWBURST_S0,
	output logic AWVALID_S0,
	input AWREADY_S0,
	
	//WRITE DATA0
	output logic [`AXI_DATA_BITS-1:0] WDATA_S0,
	output logic [`AXI_STRB_BITS-1:0] WSTRB_S0,
	output logic WLAST_S0,
	output logic WVALID_S0,
	input WREADY_S0,
	
	//WRITE RESPONSE0
	input [`AXI_IDS_BITS-1:0] BID_S0,
	input [1:0] BRESP_S0,
	input BVALID_S0,
	output logic BREADY_S0,
	
	//WRITE ADDRESS1
	output logic [`AXI_IDS_BITS-1:0] AWID_S1,
	output logic [`AXI_ADDR_BITS-1:0] AWADDR_S1,
	output logic [`AXI_LEN_BITS-1:0] AWLEN_S1,
	output logic [`AXI_SIZE_BITS-1:0] AWSIZE_S1,
	output logic [1:0] AWBURST_S1,
	output logic AWVALID_S1,
	input AWREADY_S1,
	
	//WRITE DATA1
	output logic [`AXI_DATA_BITS-1:0] WDATA_S1,
	output logic [`AXI_STRB_BITS-1:0] WSTRB_S1,
	output logic WLAST_S1,
	output logic WVALID_S1,
	input WREADY_S1,
	
	//WRITE RESPONSE1
	input [`AXI_IDS_BITS-1:0] BID_S1,
	input [1:0] BRESP_S1,
	input BVALID_S1,
	output logic BREADY_S1,
	
	//READ ADDRESS0
	output logic [`AXI_IDS_BITS-1:0] ARID_S0,
	output logic [`AXI_ADDR_BITS-1:0] ARADDR_S0,
	output logic [`AXI_LEN_BITS-1:0] ARLEN_S0,
	output logic [`AXI_SIZE_BITS-1:0] ARSIZE_S0,
	output logic [1:0] ARBURST_S0,
	output logic ARVALID_S0,
	input ARREADY_S0,
	
	//READ DATA0
	input [`AXI_IDS_BITS-1:0] RID_S0,
	input [`AXI_DATA_BITS-1:0] RDATA_S0,
	input [1:0] RRESP_S0,
	input RLAST_S0,
	input RVALID_S0,
	output logic RREADY_S0,
	
	//READ ADDRESS1
	output logic [`AXI_IDS_BITS-1:0] ARID_S1,
	output logic [`AXI_ADDR_BITS-1:0] ARADDR_S1,
	output logic [`AXI_LEN_BITS-1:0] ARLEN_S1,
	output logic [`AXI_SIZE_BITS-1:0] ARSIZE_S1,
	output logic [1:0] ARBURST_S1,
	output logic ARVALID_S1,
	input ARREADY_S1,
	
	//READ DATA1
	input [`AXI_IDS_BITS-1:0] RID_S1,
	input [`AXI_DATA_BITS-1:0] RDATA_S1,
	input [1:0] RRESP_S1,
	input RLAST_S1,
	input RVALID_S1,
	output logic RREADY_S1
	
);
    //---------- you should put your design here ----------//

	// receive
    	logic [`AXI_IDS_BITS-1:0] ARID_default;
    	logic [`AXI_ADDR_BITS-1:0] ARADDR_default;
    	logic [`AXI_LEN_BITS-1:0] ARLEN_default;
    	logic [`AXI_SIZE_BITS-1:0] ARSIZE_default;
    	logic [1:0] ARBURST_default;
    	logic ARVALID_default;
    	// send
    	logic ARREADY_default;

	// send
    	logic [`AXI_IDS_BITS-1:0] RID_default;
    	logic [`AXI_DATA_BITS-1:0] RDATA_default;
    	logic [1:0] RRESP_default;
    	logic RLAST_default;
    	logic RVALID_default;
    	// receive
    	logic RREADY_default;

	// WA receive
   	logic [`AXI_IDS_BITS-1:0] AWID_default;
   	logic [`AXI_ADDR_BITS-1:0] AWADDR_default;
   	logic [`AXI_LEN_BITS-1:0] AWLEN_default;
   	logic [`AXI_SIZE_BITS-1:0] AWSIZE_default;
   	logic [1:0] AWBURST_default;
   	logic AWVALID_default;
   	// WA send
   	logic AWREADY_default;

	// WD receive
    logic [`AXI_DATA_BITS-1:0] WDATA_default;
    logic [`AXI_STRB_BITS-1:0] WSTRB_default;
    logic WLAST_default;
    logic WVALID_default;
    // WD send
    logic WREADY_default;

	// WR send
    	logic [`AXI_IDS_BITS-1:0] BID_default;
    	logic [1:0] BRESP_default;
    	logic BVALID_default;
    	// WR receive
    	logic BREADY_default;

DefaultSlave DefaultSlave(
     .clk(ACLK),    // Clock
     .rst(ARESETn),  // Asynchronous reset active high
     // DA receive
     .ARID_default(ARID_default),
     .ARADDR_default(ARADDR_default),
     .ARLEN_default(ARLEN_default),
     .ARSIZE_default(ARSIZE_default),
     .ARBURST_default(ARBURST_default),
     .ARVALID_default(ARVALID_default),
     // DA send
     .ARREADY_default(ARREADY_default),
     // DR send
     .RID_default(RID_default),
     .RDATA_default(RDATA_default),
     .RRESP_default(RRESP_default),
     .RLAST_default(RLAST_default),
     .RVALID_default(RVALID_default),
     // DR receive
     .RREADY_default(RREADY_default),
     // WA receive
     .AWID_default(AWID_default),
     .AWADDR_default(AWADDR_default),
     .AWLEN_default(AWLEN_default),
     .AWSIZE_default(AWSIZE_default),
     .AWBURST_default(AWBURST_default),
     .AWVALID_default(AWVALID_default),
     // WA send
     .AWREADY_default(AWREADY_default),
     // WD receive
     .WDATA_default(WDATA_default),
     .WSTRB_default(WSTRB_default),
     .WLAST_default(WLAST_default),
     .WVALID_default(WVALID_default),
     // WD send
     .WREADY_default(WREADY_default),
     // WR send
     .BID_default(BID_default),
     .BRESP_default(BRESP_default),
     .BVALID_default(BVALID_default),
     // WR receive
     .BREADY_default(BREADY_default)
);



ReadAddress ReadAddress(
     .clk(ACLK),
     .rst(ARESETn),
//---------------------------master---------------------------//
     //master0 send to AXI
     .ARADDR_M0(ARADDR_M0), //data address
     .ARID_M0(ARID_M0), 
     .ARLEN_M0(ARLEN_M0),
     .ARSIZE_M0(ARSIZE_M0),
     //
     .ARBURST_M0(ARBURST_M0),
     .ARVALID_M0(ARVALID_M0),
     //M0 receive
     .ARREADY_M0(ARREADY_M0),

     //master1
     .ARADDR_M1(ARADDR_M1),
     .ARID_M1(ARID_M1),
     .ARLEN_M1(ARLEN_M1),
     .ARSIZE_M1(ARSIZE_M1),
     //
     .ARBURST_M1(ARBURST_M1),
     .ARVALID_M1(ARVALID_M1),
     //output
     .ARREADY_M1(ARREADY_M1),


//---------------------------slave---------------------------//
     //slave0 
     .ARID_S0(ARID_S0),
     .ARADDR_S0(ARADDR_S0),
     .ARLEN_S0(ARLEN_S0),
     .ARSIZE_S0(ARSIZE_S0),
     .ARVALID_S0(ARVALID_S0),
     .ARBURST_S0(ARBURST_S0),

     .ARREADY_S0(ARREADY_S0),

     //slave1 
     .ARID_S1(ARID_S1),
     .ARADDR_S1(ARADDR_S1),
     .ARLEN_S1(ARLEN_S1),
     .ARSIZE_S1(ARSIZE_S1),
     .ARVALID_S1(ARVALID_S1),
     .ARBURST_S1(ARBURST_S1),

     .ARREADY_S1(ARREADY_S1),

    //Slave default
     .ARID_default(ARID_default),
    	.ARADDR_default(ARADDR_default),
     .ARLEN_default(ARLEN_default),
    	.ARSIZE_default(ARSIZE_default),
    	.ARBURST_default(ARBURST_default),
     .ARVALID_default(ARVALID_default),
    //SlavesD send
    	.ARREADY_default(ARREADY_default)

);

ReadData Read(
     .clk(ACLK),
     .rst(ARESETn),
     //master 0 receive from AXI
     .RID_M0(RID_M0),
     .RDATA_M0(RDATA_M0),
     .RRESP_M0(RRESP_M0),
     .RLAST_M0(RLAST_M0),
     .RVALID_M0(RVALID_M0),
     //master 0 sent to slave
     .RREADY_M0(RREADY_M0),

     //master 1 receive from AXI
     .RID_M1(RID_M1),
     .RDATA_M1(RDATA_M1),
     .RRESP_M1(RRESP_M1),
     .RLAST_M1(RLAST_M1),
     .RVALID_M1(RVALID_M1),
     //master 1 sent to AXI
     .RREADY_M1(RREADY_M1),


     //SLAVE 0 sent to AXI
     .RID_S0(RID_S0),
     .RDATA_S0(RDATA_S0),
     .RRESP_S0(RRESP_S0),
     .RLAST_S0(RLAST_S0),
     .RVALID_S0(RVALID_S0),
     //master 0 sent to AXI
     .RREADY_S0(RREADY_S0),


     //SLAVE 1 
     .RID_S1(RID_S1),
     .RDATA_S1(RDATA_S1),
     .RRESP_S1(RRESP_S1),
     .RLAST_S1(RLAST_S1),
     .RVALID_S1(RVALID_S1),
     //master  sent to slave 1
     .RREADY_S1(RREADY_S1),

     //SLAVE default
     .RID_default(RID_default),
     .RDATA_default(RDATA_default),
     .RRESP_default(RRESP_default),
     .RLAST_default(RLAST_default),
     .RVALID_default(RVALID_default),
     //master  sent to slave default
     .RREADY_default(RREADY_default)

);

WriteAddress WriteAddr(
     .clk(ACLK),
     .rst(ARESETn),


     //master 1 send AXI
     .AWID_M1(AWID_M1),
     .AWADDR_M1(AWADDR_M1),
     .AWLEN_M1(AWLEN_M1),
     .AWSIZE_M1(AWSIZE_M1),
     .AWBURST_M1(AWBURST_M1),
     .AWVALID_M1(AWVALID_M1),

     //master receive
     .AWREADY_M1(AWREADY_M1),

     //slave receive from AXI
     .AWID_S0(AWID_S0),
     .AWADDR_S0(AWADDR_S0),
     .AWLEN_S0(AWLEN_S0),
     .AWSIZE_S0(AWSIZE_S0),
     .AWBURST_S0(AWBURST_S0),
     .AWVALID_S0(AWVALID_S0),
     // slave send AXI
     .AWREADY_S0(AWREADY_S0),


     .AWID_S1(AWID_S1),
     .AWADDR_S1(AWADDR_S1),
     .AWLEN_S1(AWLEN_S1),
     .AWSIZE_S1(AWSIZE_S1),
     .AWBURST_S1(AWBURST_S1),
     .AWVALID_S1(AWVALID_S1),
     // slave send
     .AWREADY_S1(AWREADY_S1),


     //slave receive firm AXI
     .AWID_default(AWID_default),
     .AWADDR_default(AWADDR_default),
     .AWLEN_default(AWLEN_default),
     .AWSIZE_default(AWSIZE_default),
     .AWBURST_default(AWBURST_default),
     .AWVALID_default(AWVALID_default),
     // slave send
     .AWREADY_default(AWREADY_default)

      
);

WriteData WriteData(
     .clk(ACLK),
     .rst(ARESETn),
     //master 0 doesn't receive data form Write data

     //master 1 to AXI

     .WDATA_M1(WDATA_M1),
     .WSTRB_M1(WSTRB_M1),
     .WLAST_M1(WLAST_M1),
     .WVALID_M1(WVALID_M1),
     // AXI to master1
     .WREADY_M1(WREADY_M1),

     //AXI to slave0
     //.WID_S0(WID_S0),
     .WDATA_S0(WDATA_S0),
     .WSTRB_S0(WSTRB_S0),
     .WLAST_S0(WLAST_S0),
     .WVALID_S0(WVALID_S0),

     .WREADY_S0(WREADY_S0),
     //AXI to slave1
     //.WID_S1(WID_S1),
     .WDATA_S1(WDATA_S1),
     .WSTRB_S1(WSTRB_S1),
     .WLAST_S1(WLAST_S1),
     .WVALID_S1(WVALID_S1),

     .WREADY_S1(WREADY_S1),

     //AXI to slave default
     //.WID_default(WID_default),
     .WDATA_default(WDATA_default),
     .WSTRB_default(WSTRB_default),
     .WLAST_default(WLAST_default),
     .WVALID_default(WVALID_default),

     .WREADY_default(WREADY_default),

     .AWVALID_S0(AWVALID_S0),
     .AWVALID_S1(AWVALID_S1),
     .AWLEN_S1(AWLEN_S1),
     /////////
     .AWVALID_default(AWVALID_default)

);

WriteRespone WriteRespone(
	.clk(ACLK),
     .rst(ARESETn),
     /*
     //master 0
     .BID_M0(BID_M0),
     .BRESP_M0(BRESP_M0),
     .BVALID_M0(BVALID_M0),
     //master 0 send
     .BREADY_M0(BREADY_M0),
     */
     //master 1
     .BID_M1(BID_M1),
     .BRESP_M1(BRESP_M1),
     .BVALID_M1(BVALID_M1),
     //master 1 send
     .BREADY_M1(BREADY_M1),

     //slave 0
     .BID_S0(BID_S0),
     .BRESP_S0(BRESP_S0),
     .BVALID_S0(BVALID_S0),
     //
     .BREADY_S0(BREADY_S0),

     //slave 0
     .BID_S1(BID_S1),
     .BRESP_S1(BRESP_S1),
     .BVALID_S1(BVALID_S1),
     //
     .BREADY_S1(BREADY_S1),

     //slave default
     .BID_default(BID_default),
     .BRESP_default(BRESP_default),
     .BVALID_default(BVALID_default),
     //
     .BREADY_default(BREADY_default)

);



endmodule
